

module cpu(

);


endmodule